magic
tech sky130A
magscale 1 2
timestamp 1687392149
<< obsli1 >>
rect 1104 2159 18860 47345
<< obsm1 >>
rect 1104 2128 19214 47376
<< obsm2 >>
rect 1582 2139 19210 47365
<< metal3 >>
rect 0 46112 800 46232
rect 19200 43392 20000 43512
rect 0 39040 800 39160
rect 0 31968 800 32088
rect 19200 31016 20000 31136
rect 0 24896 800 25016
rect 19200 18640 20000 18760
rect 0 17824 800 17944
rect 0 10752 800 10872
rect 19200 6264 20000 6384
rect 0 3680 800 3800
<< obsm3 >>
rect 800 46312 19200 47361
rect 880 46032 19200 46312
rect 800 43592 19200 46032
rect 800 43312 19120 43592
rect 800 39240 19200 43312
rect 880 38960 19200 39240
rect 800 32168 19200 38960
rect 880 31888 19200 32168
rect 800 31216 19200 31888
rect 800 30936 19120 31216
rect 800 25096 19200 30936
rect 880 24816 19200 25096
rect 800 18840 19200 24816
rect 800 18560 19120 18840
rect 800 18024 19200 18560
rect 880 17744 19200 18024
rect 800 10952 19200 17744
rect 880 10672 19200 10952
rect 800 6464 19200 10672
rect 800 6184 19120 6464
rect 800 3880 19200 6184
rect 880 3600 19200 3880
rect 800 2143 19200 3600
<< metal4 >>
rect 3163 2128 3483 47376
rect 5382 2128 5702 47376
rect 7602 2128 7922 47376
rect 9821 2128 10141 47376
rect 12041 2128 12361 47376
rect 14260 2128 14580 47376
rect 16480 2128 16800 47376
rect 18699 2128 19019 47376
<< labels >>
rlabel metal3 s 0 46112 800 46232 6 clk
port 1 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 counter[0]
port 2 nsew signal output
rlabel metal3 s 0 17824 800 17944 6 counter[1]
port 3 nsew signal output
rlabel metal3 s 0 10752 800 10872 6 counter[2]
port 4 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 counter[3]
port 5 nsew signal output
rlabel metal3 s 19200 6264 20000 6384 6 io_oeb[0]
port 6 nsew signal output
rlabel metal3 s 19200 18640 20000 18760 6 io_oeb[1]
port 7 nsew signal output
rlabel metal3 s 19200 31016 20000 31136 6 io_oeb[2]
port 8 nsew signal output
rlabel metal3 s 19200 43392 20000 43512 6 io_oeb[3]
port 9 nsew signal output
rlabel metal3 s 0 39040 800 39160 6 reset
port 10 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 up_down
port 11 nsew signal input
rlabel metal4 s 3163 2128 3483 47376 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 7602 2128 7922 47376 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 12041 2128 12361 47376 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 16480 2128 16800 47376 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 5382 2128 5702 47376 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 9821 2128 10141 47376 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 14260 2128 14580 47376 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 18699 2128 19019 47376 6 vssd1
port 13 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 696622
string GDS_FILE /home/mariam/updown_counter_openlane/openlane/mariam_updown_counter/runs/23_06_21_17_01/results/signoff/mariam_updown_counter.magic.gds
string GDS_START 144530
<< end >>

